`timescale 1ns / 1ps

module top_tb;
	parameter width=16;
	parameter N=9;
	
	reg clk;
	reg areset;
	reg signed [width-1:0] din;
	reg din_en;
	wire dout_en;
	wire [N-1:0] dout_cnt;
	wire signed [width-1:0] dout_re, dout_im;
	
	wire signed [width-1:0] dtest [(2**N-1):0];
	integer i;
	
	corefft uut (
		.clk(clk),
		.areset(areset),
		.din_en(din_en),
		.din_re(din),
		.din_im(16'd0),
		.dout_en(dout_en),
		.dout_cnt(dout_cnt),
		.dout_re(dout_re),
		.dout_im(dout_im)
	);
	
	assign dtest[0]=16'd67,
		dtest[1]=16'd64,
		dtest[2]=16'd19,
		dtest[3]=16'd13,
		dtest[4]=16'd67,
		dtest[5]=16'd108,
		dtest[6]=16'd74,
		dtest[7]=16'd3,
		dtest[8]=-16'd20,
		dtest[9]=16'd19,
		dtest[10]=16'd46,
		dtest[11]=16'd5,
		dtest[12]=-16'd57,
		dtest[13]=-16'd60,
		dtest[14]=16'd3,
		dtest[15]=16'd50,
		dtest[16]=16'd30,
		dtest[17]=-16'd8,
		dtest[18]=16'd14,
		dtest[19]=16'd88,
		dtest[20]=16'd133,
		dtest[21]=16'd102,
		dtest[22]=16'd51,
		dtest[23]=16'd57,
		dtest[24]=16'd108,
		dtest[25]=16'd120,
		dtest[26]=16'd61,
		dtest[27]=-16'd7,
		dtest[28]=-16'd8,
		dtest[29]=16'd39,
		dtest[30]=16'd51,
		dtest[31]=16'd0,
		dtest[32]=-16'd45,
		dtest[33]=-16'd17,
		dtest[34]=16'd55,
		dtest[35]=16'd85,
		dtest[36]=16'd51,
		dtest[37]=16'd22,
		dtest[38]=16'd61,
		dtest[39]=16'd128,
		dtest[40]=16'd139,
		dtest[41]=16'd82,
		dtest[42]=16'd33,
		dtest[43]=16'd50,
		dtest[44]=16'd91,
		dtest[45]=16'd75,
		dtest[46]=16'd1,
		dtest[47]=-16'd50,
		dtest[48]=-16'd26,
		dtest[49]=16'd24,
		dtest[50]=16'd20,
		dtest[51]=-16'd33,
		dtest[52]=-16'd54,
		dtest[53]=-16'd1,
		dtest[54]=16'd68,
		dtest[55]=16'd74,
		dtest[56]=16'd27,
		dtest[57]=16'd10,
		dtest[58]=16'd57,
		dtest[59]=16'd105,
		dtest[60]=16'd82,
		dtest[61]=16'd9,
		dtest[62]=-16'd29,
		dtest[63]=16'd0,
		dtest[64]=16'd29,
		dtest[65]=-16'd9,
		dtest[66]=-16'd82,
		dtest[67]=-16'd105,
		dtest[68]=-16'd57,
		dtest[69]=-16'd10,
		dtest[70]=-16'd27,
		dtest[71]=-16'd74,
		dtest[72]=-16'd68,
		dtest[73]=16'd1,
		dtest[74]=16'd54,
		dtest[75]=16'd33,
		dtest[76]=-16'd20,
		dtest[77]=-16'd24,
		dtest[78]=16'd26,
		dtest[79]=16'd50,
		dtest[80]=-16'd1,
		dtest[81]=-16'd75,
		dtest[82]=-16'd91,
		dtest[83]=-16'd50,
		dtest[84]=-16'd33,
		dtest[85]=-16'd82,
		dtest[86]=-16'd139,
		dtest[87]=-16'd128,
		dtest[88]=-16'd61,
		dtest[89]=-16'd22,
		dtest[90]=-16'd51,
		dtest[91]=-16'd85,
		dtest[92]=-16'd55,
		dtest[93]=16'd17,
		dtest[94]=16'd45,
		dtest[95]=16'd0,
		dtest[96]=-16'd51,
		dtest[97]=-16'd39,
		dtest[98]=16'd8,
		dtest[99]=16'd7,
		dtest[100]=-16'd61,
		dtest[101]=-16'd120,
		dtest[102]=-16'd108,
		dtest[103]=-16'd57,
		dtest[104]=-16'd51,
		dtest[105]=-16'd102,
		dtest[106]=-16'd133,
		dtest[107]=-16'd88,
		dtest[108]=-16'd14,
		dtest[109]=16'd8,
		dtest[110]=-16'd30,
		dtest[111]=-16'd50,
		dtest[112]=-16'd3,
		dtest[113]=16'd60,
		dtest[114]=16'd57,
		dtest[115]=-16'd5,
		dtest[116]=-16'd46,
		dtest[117]=-16'd19,
		dtest[118]=16'd20,
		dtest[119]=-16'd3,
		dtest[120]=-16'd74,
		dtest[121]=-16'd108,
		dtest[122]=-16'd67,
		dtest[123]=-16'd13,
		dtest[124]=-16'd19,
		dtest[125]=-16'd64,
		dtest[126]=-16'd67,
		dtest[127]=16'd0,
		dtest[128]=16'd67,
		dtest[129]=16'd64,
		dtest[130]=16'd19,
		dtest[131]=16'd13,
		dtest[132]=16'd67,
		dtest[133]=16'd108,
		dtest[134]=16'd74,
		dtest[135]=16'd3,
		dtest[136]=-16'd20,
		dtest[137]=16'd19,
		dtest[138]=16'd46,
		dtest[139]=16'd5,
		dtest[140]=-16'd57,
		dtest[141]=-16'd60,
		dtest[142]=16'd3,
		dtest[143]=16'd50,
		dtest[144]=16'd30,
		dtest[145]=-16'd8,
		dtest[146]=16'd14,
		dtest[147]=16'd88,
		dtest[148]=16'd133,
		dtest[149]=16'd102,
		dtest[150]=16'd51,
		dtest[151]=16'd57,
		dtest[152]=16'd108,
		dtest[153]=16'd120,
		dtest[154]=16'd61,
		dtest[155]=-16'd7,
		dtest[156]=-16'd8,
		dtest[157]=16'd39,
		dtest[158]=16'd51,
		dtest[159]=16'd0,
		dtest[160]=-16'd45,
		dtest[161]=-16'd17,
		dtest[162]=16'd55,
		dtest[163]=16'd85,
		dtest[164]=16'd51,
		dtest[165]=16'd22,
		dtest[166]=16'd61,
		dtest[167]=16'd128,
		dtest[168]=16'd139,
		dtest[169]=16'd82,
		dtest[170]=16'd33,
		dtest[171]=16'd50,
		dtest[172]=16'd91,
		dtest[173]=16'd75,
		dtest[174]=16'd1,
		dtest[175]=-16'd50,
		dtest[176]=-16'd26,
		dtest[177]=16'd24,
		dtest[178]=16'd20,
		dtest[179]=-16'd33,
		dtest[180]=-16'd54,
		dtest[181]=-16'd1,
		dtest[182]=16'd68,
		dtest[183]=16'd74,
		dtest[184]=16'd27,
		dtest[185]=16'd10,
		dtest[186]=16'd57,
		dtest[187]=16'd105,
		dtest[188]=16'd82,
		dtest[189]=16'd9,
		dtest[190]=-16'd29,
		dtest[191]=16'd0,
		dtest[192]=16'd29,
		dtest[193]=-16'd9,
		dtest[194]=-16'd82,
		dtest[195]=-16'd105,
		dtest[196]=-16'd57,
		dtest[197]=-16'd10,
		dtest[198]=-16'd27,
		dtest[199]=-16'd74,
		dtest[200]=-16'd68,
		dtest[201]=16'd1,
		dtest[202]=16'd54,
		dtest[203]=16'd33,
		dtest[204]=-16'd20,
		dtest[205]=-16'd24,
		dtest[206]=16'd26,
		dtest[207]=16'd50,
		dtest[208]=-16'd1,
		dtest[209]=-16'd75,
		dtest[210]=-16'd91,
		dtest[211]=-16'd50,
		dtest[212]=-16'd33,
		dtest[213]=-16'd82,
		dtest[214]=-16'd139,
		dtest[215]=-16'd128,
		dtest[216]=-16'd61,
		dtest[217]=-16'd22,
		dtest[218]=-16'd51,
		dtest[219]=-16'd85,
		dtest[220]=-16'd55,
		dtest[221]=16'd17,
		dtest[222]=16'd45,
		dtest[223]=16'd0,
		dtest[224]=-16'd51,
		dtest[225]=-16'd39,
		dtest[226]=16'd8,
		dtest[227]=16'd7,
		dtest[228]=-16'd61,
		dtest[229]=-16'd120,
		dtest[230]=-16'd108,
		dtest[231]=-16'd57,
		dtest[232]=-16'd51,
		dtest[233]=-16'd102,
		dtest[234]=-16'd133,
		dtest[235]=-16'd88,
		dtest[236]=-16'd14,
		dtest[237]=16'd8,
		dtest[238]=-16'd30,
		dtest[239]=-16'd50,
		dtest[240]=-16'd3,
		dtest[241]=16'd60,
		dtest[242]=16'd57,
		dtest[243]=-16'd5,
		dtest[244]=-16'd46,
		dtest[245]=-16'd19,
		dtest[246]=16'd20,
		dtest[247]=-16'd3,
		dtest[248]=-16'd74,
		dtest[249]=-16'd108,
		dtest[250]=-16'd67,
		dtest[251]=-16'd13,
		dtest[252]=-16'd19,
		dtest[253]=-16'd64,
		dtest[254]=-16'd67,
		dtest[255]=16'd0,
		dtest[256]=16'd67,
		dtest[257]=16'd64,
		dtest[258]=16'd19,
		dtest[259]=16'd13,
		dtest[260]=16'd67,
		dtest[261]=16'd108,
		dtest[262]=16'd74,
		dtest[263]=16'd3,
		dtest[264]=-16'd20,
		dtest[265]=16'd19,
		dtest[266]=16'd46,
		dtest[267]=16'd5,
		dtest[268]=-16'd57,
		dtest[269]=-16'd60,
		dtest[270]=16'd3,
		dtest[271]=16'd50,
		dtest[272]=16'd30,
		dtest[273]=-16'd8,
		dtest[274]=16'd14,
		dtest[275]=16'd88,
		dtest[276]=16'd133,
		dtest[277]=16'd102,
		dtest[278]=16'd51,
		dtest[279]=16'd57,
		dtest[280]=16'd108,
		dtest[281]=16'd120,
		dtest[282]=16'd61,
		dtest[283]=-16'd7,
		dtest[284]=-16'd8,
		dtest[285]=16'd39,
		dtest[286]=16'd51,
		dtest[287]=16'd0,
		dtest[288]=-16'd45,
		dtest[289]=-16'd17,
		dtest[290]=16'd55,
		dtest[291]=16'd85,
		dtest[292]=16'd51,
		dtest[293]=16'd22,
		dtest[294]=16'd61,
		dtest[295]=16'd128,
		dtest[296]=16'd139,
		dtest[297]=16'd82,
		dtest[298]=16'd33,
		dtest[299]=16'd50,
		dtest[300]=16'd91,
		dtest[301]=16'd75,
		dtest[302]=16'd1,
		dtest[303]=-16'd50,
		dtest[304]=-16'd26,
		dtest[305]=16'd24,
		dtest[306]=16'd20,
		dtest[307]=-16'd33,
		dtest[308]=-16'd54,
		dtest[309]=-16'd1,
		dtest[310]=16'd68,
		dtest[311]=16'd74,
		dtest[312]=16'd27,
		dtest[313]=16'd10,
		dtest[314]=16'd57,
		dtest[315]=16'd105,
		dtest[316]=16'd82,
		dtest[317]=16'd9,
		dtest[318]=-16'd29,
		dtest[319]=16'd0,
		dtest[320]=16'd29,
		dtest[321]=-16'd9,
		dtest[322]=-16'd82,
		dtest[323]=-16'd105,
		dtest[324]=-16'd57,
		dtest[325]=-16'd10,
		dtest[326]=-16'd27,
		dtest[327]=-16'd74,
		dtest[328]=-16'd68,
		dtest[329]=16'd1,
		dtest[330]=16'd54,
		dtest[331]=16'd33,
		dtest[332]=-16'd20,
		dtest[333]=-16'd24,
		dtest[334]=16'd26,
		dtest[335]=16'd50,
		dtest[336]=-16'd1,
		dtest[337]=-16'd75,
		dtest[338]=-16'd91,
		dtest[339]=-16'd50,
		dtest[340]=-16'd33,
		dtest[341]=-16'd82,
		dtest[342]=-16'd139,
		dtest[343]=-16'd128,
		dtest[344]=-16'd61,
		dtest[345]=-16'd22,
		dtest[346]=-16'd51,
		dtest[347]=-16'd85,
		dtest[348]=-16'd55,
		dtest[349]=16'd17,
		dtest[350]=16'd45,
		dtest[351]=16'd0,
		dtest[352]=-16'd51,
		dtest[353]=-16'd39,
		dtest[354]=16'd8,
		dtest[355]=16'd7,
		dtest[356]=-16'd61,
		dtest[357]=-16'd120,
		dtest[358]=-16'd108,
		dtest[359]=-16'd57,
		dtest[360]=-16'd51,
		dtest[361]=-16'd102,
		dtest[362]=-16'd133,
		dtest[363]=-16'd88,
		dtest[364]=-16'd14,
		dtest[365]=16'd8,
		dtest[366]=-16'd30,
		dtest[367]=-16'd50,
		dtest[368]=-16'd3,
		dtest[369]=16'd60,
		dtest[370]=16'd57,
		dtest[371]=-16'd5,
		dtest[372]=-16'd46,
		dtest[373]=-16'd19,
		dtest[374]=16'd20,
		dtest[375]=-16'd3,
		dtest[376]=-16'd74,
		dtest[377]=-16'd108,
		dtest[378]=-16'd67,
		dtest[379]=-16'd13,
		dtest[380]=-16'd19,
		dtest[381]=-16'd64,
		dtest[382]=-16'd67,
		dtest[383]=16'd0,
		dtest[384]=16'd67,
		dtest[385]=16'd64,
		dtest[386]=16'd19,
		dtest[387]=16'd13,
		dtest[388]=16'd67,
		dtest[389]=16'd108,
		dtest[390]=16'd74,
		dtest[391]=16'd3,
		dtest[392]=-16'd20,
		dtest[393]=16'd19,
		dtest[394]=16'd46,
		dtest[395]=16'd5,
		dtest[396]=-16'd57,
		dtest[397]=-16'd60,
		dtest[398]=16'd3,
		dtest[399]=16'd50,
		dtest[400]=16'd30,
		dtest[401]=-16'd8,
		dtest[402]=16'd14,
		dtest[403]=16'd88,
		dtest[404]=16'd133,
		dtest[405]=16'd102,
		dtest[406]=16'd51,
		dtest[407]=16'd57,
		dtest[408]=16'd108,
		dtest[409]=16'd120,
		dtest[410]=16'd61,
		dtest[411]=-16'd7,
		dtest[412]=-16'd8,
		dtest[413]=16'd39,
		dtest[414]=16'd51,
		dtest[415]=16'd0,
		dtest[416]=-16'd45,
		dtest[417]=-16'd17,
		dtest[418]=16'd55,
		dtest[419]=16'd85,
		dtest[420]=16'd51,
		dtest[421]=16'd22,
		dtest[422]=16'd61,
		dtest[423]=16'd128,
		dtest[424]=16'd139,
		dtest[425]=16'd82,
		dtest[426]=16'd33,
		dtest[427]=16'd50,
		dtest[428]=16'd91,
		dtest[429]=16'd75,
		dtest[430]=16'd1,
		dtest[431]=-16'd50,
		dtest[432]=-16'd26,
		dtest[433]=16'd24,
		dtest[434]=16'd20,
		dtest[435]=-16'd33,
		dtest[436]=-16'd54,
		dtest[437]=-16'd1,
		dtest[438]=16'd68,
		dtest[439]=16'd74,
		dtest[440]=16'd27,
		dtest[441]=16'd10,
		dtest[442]=16'd57,
		dtest[443]=16'd105,
		dtest[444]=16'd82,
		dtest[445]=16'd9,
		dtest[446]=-16'd29,
		dtest[447]=16'd0,
		dtest[448]=16'd29,
		dtest[449]=-16'd9,
		dtest[450]=-16'd82,
		dtest[451]=-16'd105,
		dtest[452]=-16'd57,
		dtest[453]=-16'd10,
		dtest[454]=-16'd27,
		dtest[455]=-16'd74,
		dtest[456]=-16'd68,
		dtest[457]=16'd1,
		dtest[458]=16'd54,
		dtest[459]=16'd33,
		dtest[460]=-16'd20,
		dtest[461]=-16'd24,
		dtest[462]=16'd26,
		dtest[463]=16'd50,
		dtest[464]=-16'd1,
		dtest[465]=-16'd75,
		dtest[466]=-16'd91,
		dtest[467]=-16'd50,
		dtest[468]=-16'd33,
		dtest[469]=-16'd82,
		dtest[470]=-16'd139,
		dtest[471]=-16'd128,
		dtest[472]=-16'd61,
		dtest[473]=-16'd22,
		dtest[474]=-16'd51,
		dtest[475]=-16'd85,
		dtest[476]=-16'd55,
		dtest[477]=16'd17,
		dtest[478]=16'd45,
		dtest[479]=16'd0,
		dtest[480]=-16'd51,
		dtest[481]=-16'd39,
		dtest[482]=16'd8,
		dtest[483]=16'd7,
		dtest[484]=-16'd61,
		dtest[485]=-16'd120,
		dtest[486]=-16'd108,
		dtest[487]=-16'd57,
		dtest[488]=-16'd51,
		dtest[489]=-16'd102,
		dtest[490]=-16'd133,
		dtest[491]=-16'd88,
		dtest[492]=-16'd14,
		dtest[493]=16'd8,
		dtest[494]=-16'd30,
		dtest[495]=-16'd50,
		dtest[496]=-16'd3,
		dtest[497]=16'd60,
		dtest[498]=16'd57,
		dtest[499]=-16'd5,
		dtest[500]=-16'd46,
		dtest[501]=-16'd19,
		dtest[502]=16'd20,
		dtest[503]=-16'd3,
		dtest[504]=-16'd74,
		dtest[505]=-16'd108,
		dtest[506]=-16'd67,
		dtest[507]=-16'd13,
		dtest[508]=-16'd19,
		dtest[509]=-16'd64,
		dtest[510]=-16'd67,
		dtest[511]=16'd0;


	initial #20000 $stop;

	initial begin
		clk <= 1;
		forever begin
			#5;
			clk <= ~clk;
		end
	end
	
	initial begin
		areset <= 1;
		#10; areset <= 0;
		#10; areset <= 1;
	end
	
	initial begin
		#21; din_en <= 1;
		for(i=0;i<(2**N-1);i=i+1) begin
			din <= dtest[i];
			#10;
		end
		din <= 16'd0;
		din_en <= 0;
	end
	
endmodule

